module vedic_8bit_multiplier(a,b,c);   
input [7:0]a;
input [7:0]b;
output [15:0]c;
wire [15:0]q0;	
wire [15:0]q1;	
wire [15:0]q2;
wire [15:0]q3;	
wire [15:0]c;
wire [7:0]temp1;
wire [11:0]temp2;
wire [11:0]temp3;
wire [11:0]temp4;
wire [7:0]q4;
wire [11:0]q5;
wire [11:0]q6;
// using 4 4x4 multipliers
vedic_4bit_multiplier z1(a[3:0],b[3:0],q0[15:0]);
vedic_4bit_multiplier z2(a[7:4],b[3:0],q1[15:0]);
vedic_4bit_multiplier z3(a[3:0],b[7:4],q2[15:0]);
vedic_4bit_multiplier z4(a[7:4],b[7:4],q3[15:0]);

// stage 1 adders 
assign temp1 ={4'b0,q0[7:4]};
adder_8bit z5(q1[7:0],temp1,q4);
assign temp2 ={4'b0,q2[7:0]};
assign temp3 ={q3[7:0],4'b0};
adder_12bit z6(temp2,temp3,q5);
assign temp4={4'b0,q4[7:0]};
// stage 2 adder
adder_12bit z7(temp4,q5,q6);
// fnal output assignment 
assign c[3:0]=q0[3:0];
assign c[15:4]=q6[11:0];



endmodule